module imem(mem_rd,data,wr_data,op1,mem_rd1,data1,wr_data1,op2,cout,clk);//module for accessing memory 16*8 
	input mem_rd,mem_rd1;//inputs
	input  [7:0]data,data1; //inputs
	input [31:0]wr_data,wr_data1; //inputs
	input clk;
	output reg cout;
	output [31:0]op1,op2;//out put
	reg [31:0]op1,op2;
	reg [31:0]address[255:0];
	reg [31:0]address1[255:0];
	//initializing address in memory
	initial
	begin
	address[0]=32'b00000000000000000000000000000000;
	address[1]=32'b00000000000000000000000000000001;
	address[2]=32'b00000000000000000000000000000010;
	address[3]=32'b00000000000000000000000000000011;
	address[4]=32'b00000000000000000000000000000100;
	address[5]=32'b00000000000000000000000000000101;
	address[6]=32'b00000000000000000000000000000110;
	address[7]=32'b00000000000000000000000000000111;
	address[8]=32'b00000000000000000000000000001000;
	address[9]=32'b00000000000000000000000000001001;
	address[10]=32'b00000000000000000000000000001010;
	address[11]=32'b00000000000000000000000000001011;
	address[12]=32'b00000000000000000000000000001100;
	address[13]=32'b00000000000000000000000000001101;
	address[14]=32'b00000000000000000000000000001110;
	address[16]=32'b00000000000000000000011101011111;
	
	address1[0]=32'b00000000000000000000000000000000;
	address1[1]=32'b00000000000000000000000000000001;
	address1[2]=32'b00000000000000000000000000000010;
	address1[3]=32'b00000000000000000000000000000011;
	address1[4]=32'b00000000000000000000000000000100;
	address1[5]=32'b00000000000000000000000000000101;
	address1[6]=32'b00000000000000000000000000000110;
	address1[7]=32'b00000000000000000000000000000111;
	address1[8]=32'b00000000000000000000000000001000;
	address1[9]=32'b00000000000000000000000000001001;
	address1[10]=32'b00000000000000000000000000001010;
	address1[11]=32'b00000000000000000000000000001011;
	address1[12]=32'b00000000000000000000000000001100;
	address1[13]=32'b00000000000000000000000000001101;
	address1[14]=32'b00000000000000000000000000001110;
	address1[16]=32'b00000000000000000000000000001111;
	address1[128]=32'b11111111111111111111111111111111;
	
	end
	always @(posedge(clk))
	begin
	  if(data[7]==1'b0)  /// instruction memory 0 to 127
	  begin
		if(!mem_rd)//memory write
		begin
		  address[data]=wr_data;
		  op1<=32'hz;
		end
		else if(mem_rd)//reading data from memory
		begin
		 op1<=address[data];
		 cout<=1'b0;
		end
		else 
		begin
		  op1<=32'hz;
		end
	  end
	
	  if(data1[7]==1'b1)/// data memory 128 to 256
	  begin
		if(!mem_rd1)//memory write
		begin
		  address1[data1]=wr_data1;
		  op2<=32'hz;
		end
		else if(mem_rd1)//reading data from memory
		begin
		 op2<=address1[data1];
		 cout<=1'b1;
		end
		else 
		begin
		  op2<=32'hz;
		end
	  end
	end
endmodule

